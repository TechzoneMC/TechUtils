// TechUtils configuration test
// Modified values follow

example1 = 112
example2 = [
    "This is",
    "stupid test"
]

example3 {
  example4 = "Yr Mum"
  example5 = "Is ugly"
}

time = "30 hours"
food = "taco"